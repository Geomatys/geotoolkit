{
 dimensions:
   lat = 4;
   lon = 2;
 variables:
   float lat(lat);
     lat:long_name = "Geodetic latitude";
     lat:units = "degrees_north";
     lat:axis = "Y";
     lat:_CoordinateAxisType = "Lat";
   float lon(lon);
     lon:long_name = "Geodetic longitude";
     lon:units = "degrees_east";
     lon:axis = "X";
     lon:_CoordinateAxisType = "Lon";
   float data(lon, lat);
 data:
lat =
  {-67.5, -22.5, 22.5, 67.5}
lon =
  {-90.0, 90.0}
data =
  {
    {0.0, 1.0, 2.0, 3.0},
    {4.0, 5.0, 6.0, 7.0}
  }
}
